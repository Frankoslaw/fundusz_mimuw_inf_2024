module cla_adder (
    input [63:0] a,
    input [63:0] b,
    input c_in,
    output c_out,
    output [63:0] sum
);
    wire [63:0] ci;

    assign ci[0] = c_in;
    assign ci[1] = (a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in));
    assign ci[2] = (a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))));
    assign ci[3] = (a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))));
    assign ci[4] = (a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))));
    assign ci[5] = (a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))));
    assign ci[6] = (a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))));
    assign ci[7] = (a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))));
    assign ci[8] = (a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))));
    assign ci[9] = (a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))));
    assign ci[10] = (a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))));
    assign ci[11] = (a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))));
    assign ci[12] = (a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))));
    assign ci[13] = (a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))));
    assign ci[14] = (a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))));
    assign ci[15] = (a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))));
    assign ci[16] = (a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))));
    assign ci[17] = (a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))));
    assign ci[18] = (a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))));
    assign ci[19] = (a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))));
    assign ci[20] = (a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))));
    assign ci[21] = (a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))));
    assign ci[22] = (a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))));
    assign ci[23] = (a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[24] = (a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[25] = (a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[26] = (a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[27] = (a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[28] = (a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[29] = (a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[30] = (a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[31] = (a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[32] = (a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[33] = (a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[34] = (a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[35] = (a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[36] = (a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[37] = (a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[38] = (a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[39] = (a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[40] = (a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[41] = (a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[42] = (a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[43] = (a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[44] = (a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[45] = (a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[46] = (a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[47] = (a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[48] = (a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[49] = (a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[50] = (a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[51] = (a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[52] = (a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[53] = (a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[54] = (a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[55] = (a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[56] = (a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[57] = (a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[58] = (a[57] & b[57]) | ((a[57] ^ b[57]) & ((a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[59] = (a[58] & b[58]) | ((a[58] ^ b[58]) & ((a[57] & b[57]) | ((a[57] ^ b[57]) & ((a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[60] = (a[59] & b[59]) | ((a[59] ^ b[59]) & ((a[58] & b[58]) | ((a[58] ^ b[58]) & ((a[57] & b[57]) | ((a[57] ^ b[57]) & ((a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[61] = (a[60] & b[60]) | ((a[60] ^ b[60]) & ((a[59] & b[59]) | ((a[59] ^ b[59]) & ((a[58] & b[58]) | ((a[58] ^ b[58]) & ((a[57] & b[57]) | ((a[57] ^ b[57]) & ((a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[62] = (a[61] & b[61]) | ((a[61] ^ b[61]) & ((a[60] & b[60]) | ((a[60] ^ b[60]) & ((a[59] & b[59]) | ((a[59] ^ b[59]) & ((a[58] & b[58]) | ((a[58] ^ b[58]) & ((a[57] & b[57]) | ((a[57] ^ b[57]) & ((a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign ci[63] = (a[62] & b[62]) | ((a[62] ^ b[62]) & ((a[61] & b[61]) | ((a[61] ^ b[61]) & ((a[60] & b[60]) | ((a[60] ^ b[60]) & ((a[59] & b[59]) | ((a[59] ^ b[59]) & ((a[58] & b[58]) | ((a[58] ^ b[58]) & ((a[57] & b[57]) | ((a[57] ^ b[57]) & ((a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    assign c_out = (a[63] & b[63]) | ((a[63] ^ b[63]) & ((a[62] & b[62]) | ((a[62] ^ b[62]) & ((a[61] & b[61]) | ((a[61] ^ b[61]) & ((a[60] & b[60]) | ((a[60] ^ b[60]) & ((a[59] & b[59]) | ((a[59] ^ b[59]) & ((a[58] & b[58]) | ((a[58] ^ b[58]) & ((a[57] & b[57]) | ((a[57] ^ b[57]) & ((a[56] & b[56]) | ((a[56] ^ b[56]) & ((a[55] & b[55]) | ((a[55] ^ b[55]) & ((a[54] & b[54]) | ((a[54] ^ b[54]) & ((a[53] & b[53]) | ((a[53] ^ b[53]) & ((a[52] & b[52]) | ((a[52] ^ b[52]) & ((a[51] & b[51]) | ((a[51] ^ b[51]) & ((a[50] & b[50]) | ((a[50] ^ b[50]) & ((a[49] & b[49]) | ((a[49] ^ b[49]) & ((a[48] & b[48]) | ((a[48] ^ b[48]) & ((a[47] & b[47]) | ((a[47] ^ b[47]) & ((a[46] & b[46]) | ((a[46] ^ b[46]) & ((a[45] & b[45]) | ((a[45] ^ b[45]) & ((a[44] & b[44]) | ((a[44] ^ b[44]) & ((a[43] & b[43]) | ((a[43] ^ b[43]) & ((a[42] & b[42]) | ((a[42] ^ b[42]) & ((a[41] & b[41]) | ((a[41] ^ b[41]) & ((a[40] & b[40]) | ((a[40] ^ b[40]) & ((a[39] & b[39]) | ((a[39] ^ b[39]) & ((a[38] & b[38]) | ((a[38] ^ b[38]) & ((a[37] & b[37]) | ((a[37] ^ b[37]) & ((a[36] & b[36]) | ((a[36] ^ b[36]) & ((a[35] & b[35]) | ((a[35] ^ b[35]) & ((a[34] & b[34]) | ((a[34] ^ b[34]) & ((a[33] & b[33]) | ((a[33] ^ b[33]) & ((a[32] & b[32]) | ((a[32] ^ b[32]) & ((a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9]) | ((a[9] ^ b[9]) & ((a[8] & b[8]) | ((a[8] ^ b[8]) & ((a[7] & b[7]) | ((a[7] ^ b[7]) & ((a[6] & b[6]) | ((a[6] ^ b[6]) & ((a[5] & b[5]) | ((a[5] ^ b[5]) & ((a[4] & b[4]) | ((a[4] ^ b[4]) & ((a[3] & b[3]) | ((a[3] ^ b[3]) & ((a[2] & b[2]) | ((a[2] ^ b[2]) & ((a[1] & b[1]) | ((a[1] ^ b[1]) & ((a[0] & b[0]) | ((a[0] ^ b[0]) & (c_in))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


    assign sum = a^b^ci;
    
endmodule